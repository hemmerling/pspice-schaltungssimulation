* D:\gruppe8\v2\transistor_acsweep_3.sch

* Schematics Version 9.1 - Web Update 1
* Thu Mar 17 10:34:42 2005



** Analysis setup **
.ac DEC 100 0.01 100000K


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "transistor_acsweep_3.net"
.INC "transistor_acsweep_3.als"


.probe


.END
